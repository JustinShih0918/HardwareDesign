module lab2_2(
    input wire clk,
    input wire rst,
    output reg [15:0] out// You can modify "reg" to "wire" if needed
);
    //Your design here

endmodule

// You can add any module you need.
// Make sure you include all modules you used in this problem.