module lab6_practice_master (
	input wire clk,
	input wire rst,
	input wire [7:0] sw, // switches
	output wire [3:0] data_out  // data (number) to slave 
);

// add your design here
endmodule

