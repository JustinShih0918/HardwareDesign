module note_gen(
    input clk, // clock from crystal
    input rst, // active high reset
    input wire [3:0] volume, 
    input [21:0] note_div_left, // div for note generation
    input [21:0] note_div_right,
    output [15:0] audio_left,
    output [15:0] audio_right
    );

    // Declare internal signals
    reg [21:0] clk_cnt_next, clk_cnt;
    reg [21:0] clk_cnt_next_2, clk_cnt_2;
    reg b_clk, b_clk_next;
    reg c_clk, c_clk_next;

    // Note frequency generation
    // clk_cnt, clk_cnt_2, b_clk, c_clk
    always @(posedge clk or posedge rst)
        if (rst == 1'b1)
            begin
                clk_cnt <= 22'd0;
                clk_cnt_2 <= 22'd0;
                b_clk <= 1'b0;
                c_clk <= 1'b0;
            end
        else
            begin
                clk_cnt <= clk_cnt_next;
                clk_cnt_2 <= clk_cnt_next_2;
                b_clk <= b_clk_next;
                c_clk <= c_clk_next;
            end
    
    // clk_cnt_next, b_clk_next
    always @*
        if (clk_cnt == note_div_left)
            begin
                clk_cnt_next = 22'd0;
                b_clk_next = ~b_clk;
            end
        else
            begin
                clk_cnt_next = clk_cnt + 1'b1;
                b_clk_next = b_clk;
            end

    // clk_cnt_next_2, c_clk_next
    always @*
        if (clk_cnt_2 == note_div_right)
            begin
                clk_cnt_next_2 = 22'd0;
                c_clk_next = ~c_clk;
            end
        else
            begin
                clk_cnt_next_2 = clk_cnt_2 + 1'b1;
                c_clk_next = c_clk;
            end

    // Assign the amplitude of the note
    // Volume is controlled here
    reg [15:0] next_high, next_low;
    reg [15:0] high, low;
    always @(posedge clk, posedge rst) begin
        if(rst) begin
            high <= 16'hDFF0;
            low <= 16'hD000;
        end
        else begin
            high <= next_high;
            low <= next_low;
        end
    end
    always @(*) begin
        if(volume == 4'b0001) begin
            next_high <= 16'hA500;
            next_low <= 16'hA000;
        end
        if(volume == 4'b0010) begin
            next_high <= 16'hDE00;
            next_low <= 16'hD500;
        end
        else if(volume == 4'b0011) begin
            next_high <= 16'hDFF0;
            next_low <= 16'hD000;
        end
        else if(volume == 4'b0100) begin
            next_high <= 16'hEE00;
            next_low <= 16'h1000;
        end
        else if(volume == 4'b0101) begin
            next_high <= 16'hE000;
            next_low <= 16'h2000;
        end
    end

    assign audio_left = (note_div_left == 22'd1) ? 16'h0000 : 
                                (b_clk == 1'b0) ? high : low;
    assign audio_right = (note_div_right == 22'd1) ? 16'h0000 : 
                                (c_clk == 1'b0) ? high : low;
endmodule