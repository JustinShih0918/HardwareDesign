`timescale 1ns/1ps
module lab2_adv_1 (
    input clk,
    input rst_n, 
    input [11:0] code, 
    output reg [3:0] out,
    output reg [7:0] raw_data,
    output reg err,
    output reg cor
);

// Output signals can be reg or wire
// add your design here
   

endmodule
