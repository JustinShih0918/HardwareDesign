module lab5_1 (
    input wire clk,
    input wire rst,
    input wire en,
    input wire dir,
    input wire vmir,
    input wire hmir,
    input wire enlarge,
    output reg [3:0] vgaRed,
    output reg [3:0] vgaGreen,
    output reg [3:0] vgaBlue,
    output reg hysnc,
    output reg vsync
);
    // add your design here

endmodule