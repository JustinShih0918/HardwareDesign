module lab6_practice_slave (
	input wire clk,
	input wire rst,
	input wire [3:0] data_in, // data (number) from master
	output wire [7:0] led // LEDs
);

// add your design here
endmodule
