module lab2_adv_2(
    input clk,
    input rst,
    input [4:0] raw_data,
    input [9:0] error_bit_input,
    output wire [9:0] received_data,
    output reg [3:0] error_index,
    output reg multiple_error
);

// Output signals can be reg or wire
// add your design here

endmodule
